module alu(
	
);



endmodule 
