module intermediateBadgeMain(

);

endmodule 